module codes

// codes color and style codes of various ansi colors and attributes.
pub const (
	black             = 30
	red               = 31
	green             = 32
	yellow            = 33
	blue              = 34
	magenta           = 35
	cyan              = 36
	white             = 37
	bright_offset     = 60
	bright_black      = 90
	bright_red        = 91
	bright_green      = 92
	bright_yellow     = 93
	bright_blue       = 94
	bright_magenta    = 95
	bright_cyan       = 96
	bright_white      = 97
	default_color     = 39
	reset             = 0
	background_offset = 10
	bold              = 1
	dim               = 2
	italic            = 3
	underline         = 4
	blinking          = 5
	inverse           = 7
	hidden            = 8
	strikethrough     = 9
)
